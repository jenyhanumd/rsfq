* RSFQ: Buffer

* assumes library/general.cir is included

.subckt buffer A B IC=.1m

    .param Ic1=1.4*IC
    .param Ib=.7*IC

    .param L=.5*Phi0/IC

    L1 A 1 L
    L2 2 B L

    xi 0 2 ibias IB=Ib

    x1 1 0 p1 cdjj IC=Ic1
    x2 2 1 p2 cdjj IC=IC

.ends buffer
